// Example macros
`define WIDTH 4
